// Code your testbench here
// or browse Examples
`timescale 1ns/1ps
`include "params_pkg.sv"

`include "axi_uvm_pkg.sv"

`include "tb.sv"
